//===========================================
// Function : The monitor module who receive
//						the data from rc6 module and 
//						then send it to the scoreboard
// FileName	: rc6_monitor.sv
// Coder    : SingularityKChen
// Edition	: edit 1
// Date     : DEC 11/2018
//===========================================